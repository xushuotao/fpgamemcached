// Copyright (c) 2013 Quanta Research Cambridge, Inc.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import MemTypes::*;
import MemServer::*;
import MMU::*;
import CtrlMux::*;
import Portal::*;
import HostInterface::*;
import ConnectalMemory::*;
import Leds::*;

// generated by tool
import BluecacheRequest::*;
import MemServerRequest::*;
import MMURequest::*;
import BluecacheIndication::*;
import MemServerIndication::*;
import MMUIndication::*;

// defined by user
import Connectable::*;
import Bluecache::*;
import DRAMCommon::*;

//import XilinxVC707DDR3::*;
`ifdef BSIM
import DDR3Sim::*;
`else
import Clocks          :: *;
import DefaultValue    :: *;
import DDR3Controller::*;
import DDR3Common::*;
//import Xilinx       :: *;
import XilinxCells ::*;
`endif
import DRAMController::*;

import AuroraCommon::*;
import ValFlashCtrlTypes::*;

//`define DDR3_VC707_1GB 29, 512, 64, 64, 8, 14, 10, 3, 1, 1, 1, 1, 1, 2

typedef enum {BluecacheIndication, BluecacheRequest, HostMemServerIndication, HostMemServerRequest, HostMMURequest, HostMMUIndication} IfcNames deriving (Eq,Bits);

interface Top_Pins;
   interface Aurora_Pins#(4) aurora_fmc1;
   interface Aurora_Clock_Pins aurora_clk_fmc1;
         
   //interface Vector#(AuroraExtQuad, Aurora_Pins#(1)) aurora_ext;
   //interface Aurora_Clock_Pins aurora_quad119;
   //interface Aurora_Clock_Pins aurora_quad117;
`ifndef BSIM
   interface DDR3_Pins_VC707_1GB pins_ddr3;
`endif
endinterface



module mkConnectalTop#(HostType host) (ConnectalTop#(PhysAddrWidth,DataBusWidth,Top_Pins,1));
   
   Clock clk250 = host.derivedClock;
   Reset rst250 = host.derivedReset;
   
   DRAMControllerIfc dramController <- mkDRAMController();
   
   `ifdef BSIM
   let ddr3_ctrl_user <- mkDDR3Simulator;
   mkConnection(dramController.ddr3_cli, ddr3_ctrl_user);

   `else 
   Clock clk200 = host.tsys_clk_200mhz_buf;
   Clock ddr_buf = clk200;
   Reset ddr3ref_rst_n <- mkAsyncResetFromCR(4, ddr_buf );
   
   DDR3_Configure ddr3_cfg = defaultValue;
   ddr3_cfg.reads_in_flight = 32;   // adjust as needed
   DDR3_Controller_VC707_1GB ddr3_ctrl <- mkDDR3Controller_VC707_2_1(ddr3_cfg, ddr_buf, clocked_by ddr_buf, reset_by ddr3ref_rst_n);
   
   Clock ddr3clk = ddr3_ctrl.user.clock;
   Reset ddr3rstn = ddr3_ctrl.user.reset_n;
   
   let ddr_cli_200Mhz <- mkDDR3ClientSync(dramController.ddr3_cli, clockOf(dramController), resetOf(dramController), ddr3clk, ddr3rstn);
   mkConnection(ddr_cli_200Mhz, ddr3_ctrl.user);
   `endif
   

   BluecacheIndicationProxy bluecacheIndicationProxy <- mkBluecacheIndicationProxy(BluecacheIndication);
   Bluecache bluecache <- mkBluecache(bluecacheIndicationProxy.ifc, clk250);
   mkConnection(bluecache.dramClient, dramController);
   BluecacheRequestWrapper bluecacheRequestWrapper <- mkBluecacheRequestWrapper(BluecacheRequest,bluecache.request);

   Vector#(1, MemReadClient#(DataBusWidth)) readClients = cons(bluecache.dmaReadClient, nil);
   Vector#(1, MemWriteClient#(DataBusWidth)) writeClients = cons(bluecache.dmaWriteClient, nil);

   MMUIndicationProxy hostMMUIndicationProxy <- mkMMUIndicationProxy(HostMMUIndication);
   MMU#(PhysAddrWidth) hostMMU <- mkMMU(0, True, hostMMUIndicationProxy.ifc);
   MMURequestWrapper hostMMURequestWrapper <- mkMMURequestWrapper(HostMMURequest, hostMMU.request);

   MemServerIndicationProxy hostMemServerIndicationProxy <- mkMemServerIndicationProxy(HostMemServerIndication);
   MemServer#(PhysAddrWidth,DataBusWidth,1) dma <- mkMemServerRW(hostMemServerIndicationProxy.ifc, readClients, writeClients, cons(hostMMU,nil));
   MemServerRequestWrapper hostMemServerRequestWrapper <- mkMemServerRequestWrapper(HostMemServerRequest, dma.request);

   Vector#(6,StdPortal) portals;
   portals[0] = hostMemServerIndicationProxy.portalIfc; 
   portals[1] = bluecacheIndicationProxy.portalIfc; 
   portals[2] = hostMemServerRequestWrapper.portalIfc;
   portals[3] = bluecacheRequestWrapper.portalIfc;
   portals[4] = hostMMURequestWrapper.portalIfc;
   portals[5] = hostMMUIndicationProxy.portalIfc;
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
   interface Top_Pins pins;
      interface Aurora_Pins aurora_fmc1 = bluecache.aurora_fmc1;
      interface Aurora_Clock_Pins aurora_clk_fmc1 = bluecache.aurora_clk_fmc1;
   
      //interface Vector#(AuroraExtQuad, Aurora_Pins#(1)) aurora_ext;
      //interface Aurora_Clock_Pins aurora_quad119;
      //interface Aurora_Clock_Pins aurora_quad117;
      `ifndef BSIM
      interface DDR3_Pins_VC707_1GB pins_ddr3 = ddr3_ctrl.ddr3;
      `endif
   endinterface


endmodule : mkConnectalTop
