import ProtocolHeader::*

