//typedef 16 NUM_STAGES;
typedef 8 NUM_STAGES;
Integer numStages = valueOf(NUM_STAGES);
