typedef 16 NUM_STAGES;
Integer numStages = valueOf(NUM_STAGES);
